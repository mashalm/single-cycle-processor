module SCProcController()